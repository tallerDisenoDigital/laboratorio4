module comparador_exponentes #(parameter bus_numero = 12, bus_exponente = 2, bus_mantisa = 8)
	(input logic[bus_numero-1:0] a,b, output logic[bus_numero-1:0] menor,mayor);
	
	
	
endmodule
